module Regfile(
  input         clock,
  input         reset,
  input         io_regWrite,
  input  [4:0]  io_rs1_s,
  input  [4:0]  io_rs2_s,
  input  [4:0]  io_rd,
  input  [31:0] io_writeData,
  output [31:0] io_rs1,
  output [31:0] io_rs2,
  output [31:0] io_regout
);
  reg [31:0] register_0; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_0;
  reg [31:0] register_1; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_1;
  reg [31:0] register_2; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_2;
  reg [31:0] register_3; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_3;
  reg [31:0] register_4; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_4;
  reg [31:0] register_5; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_5;
  reg [31:0] register_6; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_6;
  reg [31:0] register_7; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_7;
  reg [31:0] register_8; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_8;
  reg [31:0] register_9; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_9;
  reg [31:0] register_10; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_10;
  reg [31:0] register_11; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_11;
  reg [31:0] register_12; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_12;
  reg [31:0] register_13; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_13;
  reg [31:0] register_14; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_14;
  reg [31:0] register_15; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_15;
  reg [31:0] register_16; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_16;
  reg [31:0] register_17; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_17;
  reg [31:0] register_18; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_18;
  reg [31:0] register_19; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_19;
  reg [31:0] register_20; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_20;
  reg [31:0] register_21; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_21;
  reg [31:0] register_22; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_22;
  reg [31:0] register_23; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_23;
  reg [31:0] register_24; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_24;
  reg [31:0] register_25; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_25;
  reg [31:0] register_26; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_26;
  reg [31:0] register_27; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_27;
  reg [31:0] register_28; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_28;
  reg [31:0] register_29; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_29;
  reg [31:0] register_30; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_30;
  reg [31:0] register_31; // @[Regfile.scala 16:31]
  reg [31:0] _RAND_31;
  wire [31:0] _GEN_1; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_2; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_3; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_4; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_5; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_6; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_7; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_8; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_9; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_10; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_11; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_12; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_13; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_14; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_15; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_16; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_17; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_18; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_19; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_20; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_21; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_22; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_23; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_24; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_25; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_26; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_27; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_28; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_29; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_30; // @[Regfile.scala 18:16]
  wire [31:0] _GEN_33; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_34; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_35; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_36; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_37; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_38; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_39; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_40; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_41; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_42; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_43; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_44; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_45; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_46; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_47; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_48; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_49; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_50; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_51; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_52; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_53; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_54; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_55; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_56; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_57; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_58; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_59; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_60; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_61; // @[Regfile.scala 19:16]
  wire [31:0] _GEN_62; // @[Regfile.scala 19:16]
  wire  _T_2; // @[Regfile.scala 21:28]
  assign _GEN_1 = 5'h1 == io_rs1_s ? $signed(register_1) : $signed(register_0); // @[Regfile.scala 18:16]
  assign _GEN_2 = 5'h2 == io_rs1_s ? $signed(register_2) : $signed(_GEN_1); // @[Regfile.scala 18:16]
  assign _GEN_3 = 5'h3 == io_rs1_s ? $signed(register_3) : $signed(_GEN_2); // @[Regfile.scala 18:16]
  assign _GEN_4 = 5'h4 == io_rs1_s ? $signed(register_4) : $signed(_GEN_3); // @[Regfile.scala 18:16]
  assign _GEN_5 = 5'h5 == io_rs1_s ? $signed(register_5) : $signed(_GEN_4); // @[Regfile.scala 18:16]
  assign _GEN_6 = 5'h6 == io_rs1_s ? $signed(register_6) : $signed(_GEN_5); // @[Regfile.scala 18:16]
  assign _GEN_7 = 5'h7 == io_rs1_s ? $signed(register_7) : $signed(_GEN_6); // @[Regfile.scala 18:16]
  assign _GEN_8 = 5'h8 == io_rs1_s ? $signed(register_8) : $signed(_GEN_7); // @[Regfile.scala 18:16]
  assign _GEN_9 = 5'h9 == io_rs1_s ? $signed(register_9) : $signed(_GEN_8); // @[Regfile.scala 18:16]
  assign _GEN_10 = 5'ha == io_rs1_s ? $signed(register_10) : $signed(_GEN_9); // @[Regfile.scala 18:16]
  assign _GEN_11 = 5'hb == io_rs1_s ? $signed(register_11) : $signed(_GEN_10); // @[Regfile.scala 18:16]
  assign _GEN_12 = 5'hc == io_rs1_s ? $signed(register_12) : $signed(_GEN_11); // @[Regfile.scala 18:16]
  assign _GEN_13 = 5'hd == io_rs1_s ? $signed(register_13) : $signed(_GEN_12); // @[Regfile.scala 18:16]
  assign _GEN_14 = 5'he == io_rs1_s ? $signed(register_14) : $signed(_GEN_13); // @[Regfile.scala 18:16]
  assign _GEN_15 = 5'hf == io_rs1_s ? $signed(register_15) : $signed(_GEN_14); // @[Regfile.scala 18:16]
  assign _GEN_16 = 5'h10 == io_rs1_s ? $signed(register_16) : $signed(_GEN_15); // @[Regfile.scala 18:16]
  assign _GEN_17 = 5'h11 == io_rs1_s ? $signed(register_17) : $signed(_GEN_16); // @[Regfile.scala 18:16]
  assign _GEN_18 = 5'h12 == io_rs1_s ? $signed(register_18) : $signed(_GEN_17); // @[Regfile.scala 18:16]
  assign _GEN_19 = 5'h13 == io_rs1_s ? $signed(register_19) : $signed(_GEN_18); // @[Regfile.scala 18:16]
  assign _GEN_20 = 5'h14 == io_rs1_s ? $signed(register_20) : $signed(_GEN_19); // @[Regfile.scala 18:16]
  assign _GEN_21 = 5'h15 == io_rs1_s ? $signed(register_21) : $signed(_GEN_20); // @[Regfile.scala 18:16]
  assign _GEN_22 = 5'h16 == io_rs1_s ? $signed(register_22) : $signed(_GEN_21); // @[Regfile.scala 18:16]
  assign _GEN_23 = 5'h17 == io_rs1_s ? $signed(register_23) : $signed(_GEN_22); // @[Regfile.scala 18:16]
  assign _GEN_24 = 5'h18 == io_rs1_s ? $signed(register_24) : $signed(_GEN_23); // @[Regfile.scala 18:16]
  assign _GEN_25 = 5'h19 == io_rs1_s ? $signed(register_25) : $signed(_GEN_24); // @[Regfile.scala 18:16]
  assign _GEN_26 = 5'h1a == io_rs1_s ? $signed(register_26) : $signed(_GEN_25); // @[Regfile.scala 18:16]
  assign _GEN_27 = 5'h1b == io_rs1_s ? $signed(register_27) : $signed(_GEN_26); // @[Regfile.scala 18:16]
  assign _GEN_28 = 5'h1c == io_rs1_s ? $signed(register_28) : $signed(_GEN_27); // @[Regfile.scala 18:16]
  assign _GEN_29 = 5'h1d == io_rs1_s ? $signed(register_29) : $signed(_GEN_28); // @[Regfile.scala 18:16]
  assign _GEN_30 = 5'h1e == io_rs1_s ? $signed(register_30) : $signed(_GEN_29); // @[Regfile.scala 18:16]
  assign _GEN_33 = 5'h1 == io_rs2_s ? $signed(register_1) : $signed(register_0); // @[Regfile.scala 19:16]
  assign _GEN_34 = 5'h2 == io_rs2_s ? $signed(register_2) : $signed(_GEN_33); // @[Regfile.scala 19:16]
  assign _GEN_35 = 5'h3 == io_rs2_s ? $signed(register_3) : $signed(_GEN_34); // @[Regfile.scala 19:16]
  assign _GEN_36 = 5'h4 == io_rs2_s ? $signed(register_4) : $signed(_GEN_35); // @[Regfile.scala 19:16]
  assign _GEN_37 = 5'h5 == io_rs2_s ? $signed(register_5) : $signed(_GEN_36); // @[Regfile.scala 19:16]
  assign _GEN_38 = 5'h6 == io_rs2_s ? $signed(register_6) : $signed(_GEN_37); // @[Regfile.scala 19:16]
  assign _GEN_39 = 5'h7 == io_rs2_s ? $signed(register_7) : $signed(_GEN_38); // @[Regfile.scala 19:16]
  assign _GEN_40 = 5'h8 == io_rs2_s ? $signed(register_8) : $signed(_GEN_39); // @[Regfile.scala 19:16]
  assign _GEN_41 = 5'h9 == io_rs2_s ? $signed(register_9) : $signed(_GEN_40); // @[Regfile.scala 19:16]
  assign _GEN_42 = 5'ha == io_rs2_s ? $signed(register_10) : $signed(_GEN_41); // @[Regfile.scala 19:16]
  assign _GEN_43 = 5'hb == io_rs2_s ? $signed(register_11) : $signed(_GEN_42); // @[Regfile.scala 19:16]
  assign _GEN_44 = 5'hc == io_rs2_s ? $signed(register_12) : $signed(_GEN_43); // @[Regfile.scala 19:16]
  assign _GEN_45 = 5'hd == io_rs2_s ? $signed(register_13) : $signed(_GEN_44); // @[Regfile.scala 19:16]
  assign _GEN_46 = 5'he == io_rs2_s ? $signed(register_14) : $signed(_GEN_45); // @[Regfile.scala 19:16]
  assign _GEN_47 = 5'hf == io_rs2_s ? $signed(register_15) : $signed(_GEN_46); // @[Regfile.scala 19:16]
  assign _GEN_48 = 5'h10 == io_rs2_s ? $signed(register_16) : $signed(_GEN_47); // @[Regfile.scala 19:16]
  assign _GEN_49 = 5'h11 == io_rs2_s ? $signed(register_17) : $signed(_GEN_48); // @[Regfile.scala 19:16]
  assign _GEN_50 = 5'h12 == io_rs2_s ? $signed(register_18) : $signed(_GEN_49); // @[Regfile.scala 19:16]
  assign _GEN_51 = 5'h13 == io_rs2_s ? $signed(register_19) : $signed(_GEN_50); // @[Regfile.scala 19:16]
  assign _GEN_52 = 5'h14 == io_rs2_s ? $signed(register_20) : $signed(_GEN_51); // @[Regfile.scala 19:16]
  assign _GEN_53 = 5'h15 == io_rs2_s ? $signed(register_21) : $signed(_GEN_52); // @[Regfile.scala 19:16]
  assign _GEN_54 = 5'h16 == io_rs2_s ? $signed(register_22) : $signed(_GEN_53); // @[Regfile.scala 19:16]
  assign _GEN_55 = 5'h17 == io_rs2_s ? $signed(register_23) : $signed(_GEN_54); // @[Regfile.scala 19:16]
  assign _GEN_56 = 5'h18 == io_rs2_s ? $signed(register_24) : $signed(_GEN_55); // @[Regfile.scala 19:16]
  assign _GEN_57 = 5'h19 == io_rs2_s ? $signed(register_25) : $signed(_GEN_56); // @[Regfile.scala 19:16]
  assign _GEN_58 = 5'h1a == io_rs2_s ? $signed(register_26) : $signed(_GEN_57); // @[Regfile.scala 19:16]
  assign _GEN_59 = 5'h1b == io_rs2_s ? $signed(register_27) : $signed(_GEN_58); // @[Regfile.scala 19:16]
  assign _GEN_60 = 5'h1c == io_rs2_s ? $signed(register_28) : $signed(_GEN_59); // @[Regfile.scala 19:16]
  assign _GEN_61 = 5'h1d == io_rs2_s ? $signed(register_29) : $signed(_GEN_60); // @[Regfile.scala 19:16]
  assign _GEN_62 = 5'h1e == io_rs2_s ? $signed(register_30) : $signed(_GEN_61); // @[Regfile.scala 19:16]
  assign _T_2 = io_rd == 5'h0; // @[Regfile.scala 21:28]
  assign io_rs1 = 5'h1f == io_rs1_s ? $signed(register_31) : $signed(_GEN_30); // @[Regfile.scala 18:16]
  assign io_rs2 = 5'h1f == io_rs2_s ? $signed(register_31) : $signed(_GEN_62); // @[Regfile.scala 19:16]

////////////////////////////////////////////////////////////  
  assign io_regout = register_7;//                        /
////////////////////////////////////////////////////////////

`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  register_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  register_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  register_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  register_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  register_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  register_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  register_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  register_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  register_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  register_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  register_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  register_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  register_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  register_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  register_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  register_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  register_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  register_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  register_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  register_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  register_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  register_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  register_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  register_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  register_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  register_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  register_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  register_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  register_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  register_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  register_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  register_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      register_0 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          register_0 <= 32'sh0;
        end else begin
          if (5'h0 == io_rd) begin
            register_0 <= io_writeData;
          end else begin
            register_0 <= 32'sh0;
          end
        end
      end else begin
        register_0 <= 32'sh0;
      end
    end
    if (reset) begin
      register_1 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1 == io_rd) begin
            register_1 <= 32'sh0;
          end
        end else begin
          if (5'h1 == io_rd) begin
            register_1 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_2 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h2 == io_rd) begin
            register_2 <= 32'sh0;
          end
        end else begin
          if (5'h2 == io_rd) begin
            register_2 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_3 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h3 == io_rd) begin
            register_3 <= 32'sh0;
          end
        end else begin
          if (5'h3 == io_rd) begin
            register_3 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_4 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h4 == io_rd) begin
            register_4 <= 32'sh0;
          end
        end else begin
          if (5'h4 == io_rd) begin
            register_4 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_5 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h5 == io_rd) begin
            register_5 <= 32'sh0;
          end
        end else begin
          if (5'h5 == io_rd) begin
            register_5 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_6 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h6 == io_rd) begin
            register_6 <= 32'sh0;
          end
        end else begin
          if (5'h6 == io_rd) begin
            register_6 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_7 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h7 == io_rd) begin
            register_7 <= 32'sh0;
          end
        end else begin
          if (5'h7 == io_rd) begin
            register_7 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_8 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h8 == io_rd) begin
            register_8 <= 32'sh0;
          end
        end else begin
          if (5'h8 == io_rd) begin
            register_8 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_9 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h9 == io_rd) begin
            register_9 <= 32'sh0;
          end
        end else begin
          if (5'h9 == io_rd) begin
            register_9 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_10 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'ha == io_rd) begin
            register_10 <= 32'sh0;
          end
        end else begin
          if (5'ha == io_rd) begin
            register_10 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_11 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'hb == io_rd) begin
            register_11 <= 32'sh0;
          end
        end else begin
          if (5'hb == io_rd) begin
            register_11 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_12 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'hc == io_rd) begin
            register_12 <= 32'sh0;
          end
        end else begin
          if (5'hc == io_rd) begin
            register_12 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_13 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'hd == io_rd) begin
            register_13 <= 32'sh0;
          end
        end else begin
          if (5'hd == io_rd) begin
            register_13 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_14 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'he == io_rd) begin
            register_14 <= 32'sh0;
          end
        end else begin
          if (5'he == io_rd) begin
            register_14 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_15 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'hf == io_rd) begin
            register_15 <= 32'sh0;
          end
        end else begin
          if (5'hf == io_rd) begin
            register_15 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_16 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h10 == io_rd) begin
            register_16 <= 32'sh0;
          end
        end else begin
          if (5'h10 == io_rd) begin
            register_16 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_17 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h11 == io_rd) begin
            register_17 <= 32'sh0;
          end
        end else begin
          if (5'h11 == io_rd) begin
            register_17 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_18 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h12 == io_rd) begin
            register_18 <= 32'sh0;
          end
        end else begin
          if (5'h12 == io_rd) begin
            register_18 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_19 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h13 == io_rd) begin
            register_19 <= 32'sh0;
          end
        end else begin
          if (5'h13 == io_rd) begin
            register_19 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_20 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h14 == io_rd) begin
            register_20 <= 32'sh0;
          end
        end else begin
          if (5'h14 == io_rd) begin
            register_20 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_21 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h15 == io_rd) begin
            register_21 <= 32'sh0;
          end
        end else begin
          if (5'h15 == io_rd) begin
            register_21 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_22 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h16 == io_rd) begin
            register_22 <= 32'sh0;
          end
        end else begin
          if (5'h16 == io_rd) begin
            register_22 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_23 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h17 == io_rd) begin
            register_23 <= 32'sh0;
          end
        end else begin
          if (5'h17 == io_rd) begin
            register_23 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_24 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h18 == io_rd) begin
            register_24 <= 32'sh0;
          end
        end else begin
          if (5'h18 == io_rd) begin
            register_24 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_25 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h19 == io_rd) begin
            register_25 <= 32'sh0;
          end
        end else begin
          if (5'h19 == io_rd) begin
            register_25 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_26 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1a == io_rd) begin
            register_26 <= 32'sh0;
          end
        end else begin
          if (5'h1a == io_rd) begin
            register_26 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_27 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1b == io_rd) begin
            register_27 <= 32'sh0;
          end
        end else begin
          if (5'h1b == io_rd) begin
            register_27 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_28 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1c == io_rd) begin
            register_28 <= 32'sh0;
          end
        end else begin
          if (5'h1c == io_rd) begin
            register_28 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_29 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1d == io_rd) begin
            register_29 <= 32'sh0;
          end
        end else begin
          if (5'h1d == io_rd) begin
            register_29 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_30 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1e == io_rd) begin
            register_30 <= 32'sh0;
          end
        end else begin
          if (5'h1e == io_rd) begin
            register_30 <= io_writeData;
          end
        end
      end
    end
    if (reset) begin
      register_31 <= 32'sh0;
    end else begin
      if (io_regWrite) begin
        if (_T_2) begin
          if (5'h1f == io_rd) begin
            register_31 <= 32'sh0;
          end
        end else begin
          if (5'h1f == io_rd) begin
            register_31 <= io_writeData;
          end
        end
      end
    end
  end
endmodule